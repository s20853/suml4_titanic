���9      �sklearn.ensemble._forest��RandomForestClassifier���)��}�(�	estimator��sklearn.tree._classes��DecisionTreeClassifier���)��}�(�	criterion��gini��splitter��best��	max_depth�N�min_samples_split�K�min_samples_leaf�K�min_weight_fraction_leaf�G        �max_features�N�max_leaf_nodes�N�random_state�N�min_impurity_decrease�G        �class_weight�N�	ccp_alpha�G        �_sklearn_version��1.2.2�ub�n_estimators�K
�estimator_params�(hhhhhhhhhht��base_estimator��
deprecated��	bootstrap���	oob_score���n_jobs�NhK:�verbose�K �
warm_start��hN�max_samples�NhhhKhKhKhG        h�sqrt�hNhG        hG        �feature_names_in_��numpy.core.multiarray��_reconstruct����numpy��ndarray���K ��Cb���R�(KK��h+�dtype����O8�����R�(K�|�NNNJ����J����K?t�b�]�(�Pclass��Sex��Age��SibSp��Parch��Fare��Embarked�et�b�n_features_in_�K�
n_outputs_�K�classes_�h*h-K ��h/��R�(KK��h4�i8�����R�(K�<�NNNJ����J����K t�b�C               �t�b�
n_classes_�K�
estimator_�h	�estimators_�]�(h)��}�(hhhhhKhKhKhG        hh&hNhJ#�w]hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h4�f8�����R�(KhMNNNJ����J����K t�b�C              �?�t�bhQh(�scalar���hLC       ���R��max_features_�K�tree_��sklearn.tree._tree��Tree���Kh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hK�
node_count�K�nodes�h*h-K ��h/��R�(KK��h4�V56�����R�(Kh8N(�
left_child��right_child��feature��	threshold��impurity��n_node_samples��weighted_n_node_samples�t�}�(h}h4�i8�����R�(KhMNNNJ����J����K t�bK ��h~h�K��hh�K��h�h]K��h�h]K ��h�h�K(��h�h]K0��uK8KKt�b�BH                          �TL@�'�H��?�           8�@                        ��Y"@8&f.)�?�           �@                          �;@b:�&���?�             o@������������������������       ��/�L���?>            @W@������������������������       �0����a�?c            �c@                           �?��n�u�?�            �v@������������������������       ��b�{�?]            `a@������������������������       �*�8�4�?�            �k@	                        @3[Q@��Q��?B             Y@
                          �M@�KM�]�?             3@������������������������       �        
             1@������������������������       �                      @                          �E@�5��?7            @T@������������������������       �.Lj���?/             Q@������������������������       ��θ�?             *@�t�b�values�h*h-K ��h/��R�(KKKK��h]�C�     p}@      n@     @{@     �e@     �i@     �F@     �P@      :@      a@      3@      m@     @`@      I@     @V@     �f@     �D@     �A@     @P@       @      1@              1@       @             �@@      H@      7@     �F@      $@      @�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ [UhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                             �?��ϙLq�?�           8�@                          �?@��F3��?�             o@                           @�7�?s            �g@������������������������       ��|G7�?e            �d@������������������������       ����|���?             6@                            @�r����?,             N@������������������������       � ��WV�?%             J@������������������������       �      �?              @	                           +@4�^���?           �|@
                           �?�q�q�?             ;@������������������������       ��q�q�?             @������������������������       ����N8�?             5@                           �?�r����?	           0{@������������������������       �r٣����?%            �P@������������������������       �����X��?�            w@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�     �|@     �o@     �Q@     `f@      O@     �_@      H@     �]@      ,@       @       @      J@       @      I@      @       @      x@      S@      "@      2@      @       @      @      0@     �w@      M@      I@      0@     pt@      E@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ;�shG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                              @�4�O��?�           8�@                           �?�L�����?�            �t@                           �?��&�=��?�            �j@������������������������       �����1�?+            @R@������������������������       �qb����?V            �a@                          kp@��5Վ3�?S            �]@������������������������       �Dc}h��?O             \@������������������������       �����X�?             @	                        pff@=87��?�            �w@
                        �|Y;@�h����?%             L@������������������������       ��LQ�1	�?             7@������������������������       �                    �@@                           @���z��?�             t@������������������������       �     ��?             0@������������������������       ��K�)���?�             s@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�     �{@     �p@      c@     �f@     @\@     @Y@      @     �P@     �Z@     �A@     �C@      T@      A@     �S@      @       @     pr@     �T@     �J@      @      4@      @     �@@             @n@      T@      @      "@     `m@     �Q@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ\0dhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                             �?n��"�)�?�           8�@                          �;@�)z� ��?X            `a@                           @ s�n_Y�?             J@������������������������       �                     @������������������������       ���Hg���?            �F@                           �?f?8���?9            �U@������������������������       �`Jj��?             ?@������������������������       �d}h���?#             L@	                           @��O�A�?h           ��@
                            @�0�.w�?Z            �@������������������������       ��f���?�             o@������������������������       ����C�?�            �r@                           �?�8��8��?             8@������������������������       �z�G�z�?             $@������������������������       �        
             ,@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�     �y@     �r@     �L@     �T@      &@     �D@              @      &@      A@      G@     �D@       @      =@      F@      (@     @v@      k@     �t@     �j@     �[@     @a@     �k@      S@      6@       @       @       @      ,@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ���~hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                             �?"��p�?�           8�@                            @ڤ���?�            `n@                           @5�wAd�?V            �`@������������������������       ��q�q�?             @������������������������       ��z�N��?T            ``@                           @�A�|O��?C            @[@������������������������       ��[�IJ�?;            �W@������������������������       �                     .@	                            �?�i� ���?           @}@
                           2@���!x��?;            @Y@������������������������       �                     "@������������������������       � �&�T�?7             W@                           �?pH?�U��?�            �v@������������������������       ����c���?�            �s@������������������������       ���N`.�?$            �K@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�      {@     Pq@      N@     �f@      @      `@       @      �?      @      `@     �K@      K@      D@      K@      .@             `w@     �W@     �P@      A@              "@     �P@      9@     0s@      N@     �p@      E@     �B@      2@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�kfvhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtK	huh*h-K ��h/��R�(KK	��h|�B�                            @M@��l�Qf�?�           8�@                           �?�ت��?�           x�@                        `f�$@*O���?+           @}@������������������������       � �y63��?�            �n@������������������������       ��2�QZ��?�            �k@                           �?rl[غ��?�            `k@������������������������       �ڷv���?I            �\@������������������������       �҆�s��?C             Z@������������������������       �                     8@�t�bh�h*h-K ��h/��R�(KK	KK��h]�C�     0{@     @q@     �y@     @q@     �r@      e@     �h@     �G@     @Y@     �^@      \@     �Z@     �E@      R@     @Q@     �A@      8@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ��[hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                              @|��;;��?�           8�@                           �?�'�G�V�?�            �s@                            �?�Y�R_�?+            �Q@������������������������       ��4��?'            @P@������������������������       �                     @                          �(@�r�����?�            @n@������������������������       ��t����?             A@������������������������       �z0��k��?x             j@	                           �?�:,&�e�?�            �x@
                        �|>@z0��k��??             Z@������������������������       �lG:<�?:            @X@������������������������       �                     @                           @R�?�*�?�            `r@������������������������       �꒹H���?�            �q@������������������������       �        	             ,@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�     �z@     �q@     �`@     `f@      6@     �H@      6@     �E@              @      \@     @`@      >@      @     �T@     �_@     �r@     �Y@     �O@     �D@      L@     �D@      @              m@     �N@     `k@     �N@      ,@        �t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�nwhG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                           xWI@"��p�?�           8�@                           �?�A����?�           ��@                           �?���i!��?z            `f@������������������������       � \� ���?'            �H@������������������������       �6�z���?S            @`@                           *@��0���?           �y@������������������������       ��P�*�?             ?@������������������������       �0%���?�?�            �w@	                           �?^;|��?Q            �]@
                           �?L紂P�?"            �I@������������������������       �                     @@������������������������       �p�ݯ��?             3@                           �?ҳ�wY;�?/             Q@������������������������       ��ݜ�?            �C@������������������������       �J�8���?             =@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�      {@     Pq@     0y@     �g@     @P@     �\@      (@     �B@     �J@     @S@      u@     �R@      *@      2@     Pt@     �L@      ?@      V@      @      F@              @@      @      (@      8@      F@      @      A@      3@      $@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ��^hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                             �?e�L��?�           8�@                           @�)V���?�            �p@                          �?@
ҵR�?�            Pp@������������������������       �Zw6G���?o            `f@������������������������       �������?0            �T@                          @C@r�q��?             @������������������������       �      �?              @������������������������       �                     @	                        �?�@�Y�?�(�?           �{@
                          �;@DgV`�?T            ``@������������������������       ��8��8��?!             H@������������������������       � Df@��?3            �T@                           �?\fc9�?�            �s@������������������������       �     ��?#             P@������������������������       ��w>�
��?�             o@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�     �{@     �p@     �R@      h@     �Q@     �g@      O@     @]@       @     �R@      @      �?      �?      �?      @              w@      S@     @_@      @      F@      @     @T@       @     `n@     �Q@      E@      6@      i@      H@�t�bubhhubh)��}�(hhhhhKhKhKhG        hh&hNhJ�x�	hG        hNhG        hCKhDKhEh*h-K ��h/��R�(KK��h]�C              �?�t�bhQhbhLC       ���R�hfKhghjKh*h-K ��h/��R�(KK��hL�C       �t�bK��R�}�(hKhtKhuh*h-K ��h/��R�(KK��h|�BH                          `f�$@^����[�?�           8�@                           �?�~�4_��?�            �p@                           -@���|���?#            �K@������������������������       �؇���X�?             @������������������������       ��q�q�?              H@                            @�KM�]�?�             j@������������������������       �                     $@������������������������       �$%��5,�?�            �h@	                            @@s�
��?           �{@
                           �?�D�	9�?�            @s@������������������������       ���ZE��?�            �j@������������������������       �r�q��?7             X@                          �*@�^�!<�?V            `a@������������������������       �                      @������������������������       ��nU���?P            ``@�t�bh�h*h-K ��h/��R�(KKKK��h]�C�     @{@     0q@     �i@     �L@      4@     �A@      @      �?      ,@      A@     `g@      6@      $@              f@      6@     �l@     @k@     @`@     @f@     @Z@     �Z@      9@     �Q@     �X@      D@               @     �X@      @@�t�bubhhubehhub.